module MixColumns(

);


endmodule
