module Decrypt(
input [127:0] SecretKey,
input [127:0] PlainText,
input clk,
output [127:0] CipherText
);
//order
InvShiftRows()
InvSubBytes()
InvMixColumns

endmodule
