module load_matrices();
// TODO(arianaolson419): Implement!
endmodule