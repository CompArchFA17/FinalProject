module SBoxLookup(

input num,
output outnum 

); 

reg out;
wire [1:0] in;


always @(in)
case(in)
		// source fopr s box is http://www.samiam.org/s-box.html 
	8'b000 		: out = 01100011; //63		// did Logan count in binary correctly? 
	8'b001 		: out = 01111100; //7c				// the world may never know 
	8'b010 		: out = 01110111; //77 
	8'b011 		: out = 01111011; //7b
	8'b100 		: out = 11110010; //f2
	8'b101 		: out = 01101011; //6b
	8'b110 		: out = 01101111; //6f
	8'b111 		: out = 11000101; //c5
	8'b1000 	: out = 00110000; //30
	8'b1001 	: out = 00000001; //01
	8'b1010 	: out = 01100111; //67
	8'b1011 	: out = 00101011; //2b
	8'b1100 	: out = 11111110; //fe
	8'b1101 	: out = 11010111; //d7
	8'b1110 	: out = 10101011; //ab
	8'b1111 	: out = 01110110; //76     // end of first row 
	
	8'b10000 	: out = ; // ca
	8'b10001 	: out = ; // 82
	8'b10010 	: out = ; // c9
	8'b10011 	: out = ; // 7d
	8'b10100 	: out = ; // fa
	8'b10101 	: out = ; // 59
	8'b10110 	: out = ; // 47
	8'b10111 	: out = ; // f0
	8'b11000 	: out = ; // ad
	8'b11001 	: out = ; // d4
	8'b11010 	: out = ; // a2
	8'b11011 	: out = ; // af
	8'b11100 	: out = ; // 9c
	8'b11101 	: out = ; // a4
	8'b11110 	: out = ; // 72
	8'b11111 	: out = ; // c0		// end of second row 
	
	
	8'b100001 	: out = ; // b7
	8'b100010 	: out = ; // fd
	8'b100011 	: out = ; // 93
	8'b100100 	: out = ; // 26
	8'b100101 	: out = ; // 36
	8'b100110 	: out = ; // 3f
	8'b100111 	: out = ; // f7
	8'b101000 	: out = ; // cc
	8'b101001 	: out = ; // 34
	8'b101010 	: out = ; // a5
	8'b101011 	: out = ; // e5
	8'b101100 	: out = ; // f1
	8'b101101 	: out = ; // 71
	8'b101110 	: out = ; // d8
	8'b101111 	: out = ; // 31
	8'b110000 	: out = ; // 15		// end of third row 
	
	
	8'b110001 	: out = ; // 04
	8'b110010 	: out = ; // c7
	8'b110011 	: out = ; // 23
	8'b110100 	: out = ; // c3
	8'b110101 	: out = ; // 18
	8'b110110 	: out = ; // 96
	8'b110111 	: out = ; // 05
	8'b111000 	: out = ; // 9a
	8'b111001 	: out = ; // 07
	8'b111010 	: out = ; // 12
	8'b111011 	: out = ; // 80
	8'b111100 	: out = ; // e2
	8'b111101 	: out = ; // eb
	8'b111110 	: out = ; // 27
	8'b111111 	: out = ; // b2
	8'b1000000 	: out = ; // 75// 4th row
	
	
	8'b1000001 	: out = ; // 09
	8'b1000010 	: out = ; // 83
	8'b1000011 	: out = ; // 2c
	8'b1000100 	: out = ; // 1a
	8'b1000101 	: out = ; // 1b
	8'b1000110 	: out = ; // 6e
	8'b1000111 	: out = ; // 5a
	8'b1001000 	: out = ; // a0
	8'b1001001 	: out = ; // 52
	8'b1001010 	: out = ; // 3b
	8'b1001011 	: out = ; // d6
	8'b1001100 	: out = ; // b3
	8'b1001101 	: out = ; // 29
	8'b1001110 	: out = ; // e3
	8'b1001111 	: out = ; // 2f
	8'b1010000 	: out = ; // 84		/5th row
	
	
	8'b1010001 	: out = ; // 53
	8'b1010010 	: out = ; // d1
	8'b1010011 	: out = ; // 00
	8'b1010100 	: out = ; // ed
	8'b1010101 	: out = ; // 20
	8'b1010110 	: out = ; // fc
	8'b1010111 	: out = ; // b1
	8'b1011000 	: out = ; // 5b
	8'b1011001 	: out = ; // 6a
	8'b1011010 	: out = ; // cb
	8'b1011011 	: out = ; // be
	8'b1011100 	: out = ; // 39
	8'b1011101 	: out = ; // 4a
	8'b1011110 	: out = ; // 4c
	8'b1011111 	: out = ; // 58
	8'b1100000 	: out = ; // cf		// 6th row 
	
	
	8'b1100001 	: out = ; // d0
	8'b1100010 	: out = ; // ef
	8'b1100011 	: out = ; // aa
	8'b1100100 	: out = ; // fb
	8'b1100101 	: out = ; // 43
	8'b1100110 	: out = ; // 4d
	8'b1100111 	: out = ; // 33
	8'b1101000 	: out = ; // 85
	8'b1101001 	: out = ; // 45
	8'b1101010 	: out = ; // f9
	8'b1101011 	: out = ; // 02
	8'b1101100 	: out = ; // 7f
	8'b1101101 	: out = ; // 50
	8'b1101110 	: out = ; // 3c
	8'b1101111 	: out = ; // 9f
	8'b1110000 	: out = ; // a8		/7th row 
	
	
	8'b1000000 	: out = ; // 51
	8'b1000000 	: out = ; // a3
	8'b1000000 	: out = ; // 40
	8'b1000000 	: out = ; // 8f
	8'b1000000 	: out = ; // 92
	8'b1000000 	: out = ; // 9d
	8'b1000000 	: out = ; // 38
	8'b1000000 	: out = ; // f5
	8'b1000000 	: out = ; // bc
	8'b1000000 	: out = ; // b6
	8'b1000000 	: out = ; // da
	8'b1000000 	: out = ; // 21
	8'b1000000 	: out = ; // 10
	8'b1000000 	: out = ; // ff
	8'b1000000 	: out = ; // f3
	8'b1000000 	: out = ; // d2		//8th row 
	
	
	8'b1000000 	: out = ; // cd
	8'b1000000 	: out = ; // 0c
	8'b1000000 	: out = ; // 13
	8'b1000000 	: out = ; // ec
	8'b1000000 	: out = ; // 5f
	8'b1000000 	: out = ; // 97
	8'b1000000 	: out = ; // 44
	8'b1000000 	: out = ; // 17
	8'b1000000 	: out = ; // c4
	8'b1000000 	: out = ; // a7
	8'b1000000 	: out = ; // 7e
	8'b1000000 	: out = ; // 3d
	8'b1000000 	: out = ; // 64
	8'b1000000 	: out = ; // 5d
	8'b1000000 	: out = ; // 19
	8'b1000000 	: out = ; // 73		// 9th row 
	
	
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	8'b1000000 	: out = ; // 
	
	

	
	
	
	
	 
		
	



endcase



endmodule 
