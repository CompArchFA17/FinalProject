module ShiftRows(

);

endmodule
