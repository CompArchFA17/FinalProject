module ShiftRows(

);



endmodule
